//Make your struct here


class alu_data;
        //Initialize your struct here


        // Class methods(tasks) go here


        // Constraints


endclass: alu_data

